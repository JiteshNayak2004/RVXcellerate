module top(input logic clk, reset,
			  output logic [31:0] writedata, dataadr,
			  output logic 		 memwrite);
			  
	logic [31:0] pc, instr, readdata;
	
	risc r1(clk, reset, pc, instr, memwrite, dataadr,
			  writedata, readdata);
	
	imem i1(pc[7:2], instr);
	
	dmem d1(clk, memwrite, dataadr, writedata, readdata);

endmodule 